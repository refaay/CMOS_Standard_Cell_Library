*** SPICE deck for cell osc5{sch} from library Project1
*** Created on Sun Apr 01, 2018 22:23:49
*** Last revised on Sun Apr 01, 2018 22:43:14
*** Written on Sun Apr 01, 2018 22:43:25 by Electric VLSI Design System, version 9.07
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

*** SUBCIRCUIT Project1__inv_1 FROM CELL Project1:inv_1{sch}
.SUBCKT Project1__inv_1 in out
** GLOBAL gnd
** GLOBAL vdd
Mnmos@1 out in gnd gnd N L=0.2U W=0.3U
Mpmos@0 vdd in out vdd P L=0.2U W=0.6U
.ENDS Project1__inv_1

.global gnd vdd

*** TOP LEVEL CELL: Project1:osc5{sch}
Xinv_1@0 out net@0 Project1__inv_1
Xinv_1@1 net@0 net@1 Project1__inv_1
Xinv_1@2 net@1 net@2 Project1__inv_1
Xinv_1@3 net@2 net@3 Project1__inv_1
Xinv_1@4 net@3 out Project1__inv_1
Xinv_1@6 inv_1@6_in inv_1@6_out Project1__inv_1

* Spice Code nodes in cell cell 'Project1:osc5{sch}'
vsupply vdd 0 3.3v
vgnd gnd 0 0v
.include C:\Electric\scmos18.txt
.tran 0.01ns 5ns
* Dummy control block for SPICE 3
.control
.endc
.END
